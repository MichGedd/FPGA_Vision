module system(input a, output x);
	assign x = a;
endmodule
