module system(input [7:0] a, output [7:0] x);
	assign x = a;
endmodule
